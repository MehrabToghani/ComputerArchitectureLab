module DFlipFlop;
	initial begin
		$display("Init");
	end
endmodule
